`timescale 1ns / 1ps

module CPU_RV32I (
    input  logic        clk,
    input  logic        reset,
    input  logic [31:0] instrCode,
    output logic [31:0] instrMemAddr,
    output logic        busWe,
    output logic [31:0] busAddr,
    output logic [31:0] busWData,
    input  logic [31:0] busRData
);

    logic       regFileWe;
    logic [3:0] aluControl;
    logic       aluSrcMuxSel;
    logic [1:0] RFWDSrcMuxSel;
    logic       branch;
    logic       RD1MuxSel;
    logic       jump;

    ControlUnit U_ControlUnit (.*);
    DataPath U_DataPath (.*);
endmodule
