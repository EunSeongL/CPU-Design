// Register File
`define RF_PATH   U_MCU.U_CPU_RV32I.U_DataPath.U_RegFile

// Instruction Memory
`define INSTR_PATH U_MCU.U_ROM

// Data Memory
`define RAM_PATH  U_MCU.U_RAM

