`define  ADD      4'b0000    //  ADD
`define  SUB      4'b1000    //  SUB
`define  SLL      4'b0001    //  SLL
`define  SRL      4'b0101    //  SRL
`define  SRA      4'b1101    //  SRA
`define  SLT      4'b0010    //  SLT
`define SLTU      4'b0011    // SLTU
`define  XOR      4'b0100    //  XOR
`define   OR      4'b0110    //   OR
`define  AND      4'b0111    //  AND

`define OP_TYPE_R 7'b0110011 // R-Type
`define OP_TYPE_S 7'b0100011 // S-Type
`define OP_TYPE_L 7'b0000011 // L-Type
`define OP_TYPE_I 7'b0010011 // I-Type

